/*
 *Author: vani2620
 *Date created: 24012025
*/

// verilog_lint: waive-start macro-name-style
// verilog_lint: waive-start parameter-name-style

`ifndef alpharetz_uart_params
`define alpharetz_uart_params
parameter int UART_DATA_WIDTH = 8;
parameter shortint UART_CLK_RATIO = 16;
`endif
